`timescale 1ns / 1ps
module main(
    input clk,
    input reset,
    input Start_K_G,
    output end_K_G
    );
endmodule

`timescale 1ns / 1ps
module matrix_inversion(

    );
endmodule
